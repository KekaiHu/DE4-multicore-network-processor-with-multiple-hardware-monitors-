//
// Designed by Qiang Wu
//	16K bytes, 32bit interface

`timescale 1ns/1ps


module localram(clk, addr, data_in, data_out, we, en, reset);
input clk;
input [13:2] addr;
input [31:0] data_in;
output [31:0] data_out;
input [3:0] we;
input en;
input reset;


RAMB16_S4 localram0(
	.DO     (data_out[3:0]),
	.ADDR   (addr[13:2]),
	.CLK    (clk),
	.DI     (data_in[3:0]),
	.EN     (en),
	.SSR    (reset),
	.WE     (we[0])
);
defparam localram0.INIT_00 = 256'hCA40C840C8404001C840C840C840CA40C840C840400409014DA0804000000203;
defparam localram0.INIT_01 = 256'h002000000C0002044200000400C1000040C81480884114808010C840C840C840;
defparam localram0.INIT_02 = 256'h41060C1208C2001C0008F001C0008C0704810C0000CC20000080CF0000040030;
defparam localram0.INIT_03 = 256'h00100004FF0000C00F000080854880000D040750001000C00808508880008008;
defparam localram0.INIT_04 = 256'h0000000001000000050010040F000000040040F410407AF4420000000000C005;
defparam localram0.INIT_05 = 256'h4101041041410041041441004104104104444444400000000000000000000000;
defparam localram0.INIT_06 = 256'h0000041041041041041041044101041041410404104141004104104104104104;
defparam localram0.INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;


RAMB16_S4 localram1(
	.DO     (data_out[7:4]),
	.ADDR   (addr[13:2]),
	.CLK    (clk),
	.DI     (data_in[7:4]),
	.EN     (en),
	.SSR    (reset),
	.WE     (we[0])
);
defparam localram1.INIT_00 = 256'h3333222211110005666655554444333322221111009105000F20F00000000100;
defparam localram1.INIT_01 = 256'h0000000001000C011000000100F00000013323C0000220F00007666655554444;
defparam localram1.INIT_02 = 256'h20010020010000258010F0025801000D121201220021000000202F00000200B0;
defparam localram1.INIT_03 = 256'h00200002FF0000100F0000202202200000020C60110010D00202202020000000;
defparam localram1.INIT_04 = 256'h0000000600000020020020000F00000200000010000002F00000000200001002;
defparam localram1.INIT_05 = 256'h0010100100001100100000110010010010000000000000000000000000000000;
defparam localram1.INIT_06 = 256'h0000100100100100100100100010100100001010010000110010010010010010;
defparam localram1.INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;


RAMB16_S4 localram2(
	.DO     (data_out[11:8]),
	.ADDR   (addr[13:2]),
	.CLK    (clk),
	.DI     (data_in[11:8]),
	.EN     (en),
	.SSR    (reset),
	.WE     (we[1])
);
defparam localram2.INIT_00 = 256'h000000000000000000000000000000000000000000F000000F80F08080800000;
defparam localram2.INIT_01 = 256'h002F0000000000800400000000F00F08000000F0000800F00000000000000000;
defparam localram2.INIT_02 = 256'h00000082000200050000000050000000000000004000400000000F0000000000;
defparam localram2.INIT_03 = 256'h008200000F0000000F0000000000000000000F00000000000000000000000400;
defparam localram2.INIT_04 = 256'h0000000000800000000084000F00000000100010100000E00400000000000000;
defparam localram2.INIT_05 = 256'h1118765432111DCBA987111321FEDC1111111111100000000000000000000000;
defparam localram2.INIT_06 = 256'h0000BA98765432111DCBA987111321FEDC1118765432111DCBA987111321FEDC;
defparam localram2.INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;


RAMB16_S4 localram3(
	.DO     (data_out[15:12]),
	.ADDR   (addr[13:2]),
	.CLK    (clk),
	.DI     (data_in[15:12]),
	.EN     (en),
	.SSR    (reset),
	.WE     (we[1])
);
defparam localram3.INIT_00 = 256'h000000000000000000000000000000000000000000F000600F10101010100000;
defparam localram3.INIT_01 = 256'h001F0000001000000100000010F001010000F0F0000EF0F60700000000000000;
defparam localram3.INIT_02 = 256'h00000011000100102000000102000000000100001000100000010F0000001000;
defparam localram3.INIT_03 = 256'h001100010F0000010F0000010100000100000F00000000000010100000010100;
defparam localram3.INIT_04 = 256'h0000000000100001010011000F00000010000000000001F00100000010000101;
defparam localram3.INIT_05 = 256'h0002222222000111111100011100000000000000000000000000000000000000;
defparam localram3.INIT_06 = 256'h0000666666666600055555550005554444000444444400033333330003332222;
defparam localram3.INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;


RAMB16_S4 localram4(
	.DO     (data_out[19:16]),
	.ADDR   (addr[13:2]),
	.CLK    (clk),
	.DI     (data_in[19:16]),
	.EN     (en),
	.SSR    (reset),
	.WE     (we[2])
);
defparam localram4.INIT_00 = 256'hEDCBA98765432100F9876543210FEDCBA987654321D000884050DD5544CC0000;
defparam localram4.INIT_01 = 256'h2222022022200223220220222022320200540ED00DE00EDA0BADF9876543210F;
defparam localram4.INIT_02 = 256'h2202020202220222232220222232000000220232202220220222220220222000;
defparam localram4.INIT_03 = 256'h0202022222320222220220232223202200020020222020020232302320222202;
defparam localram4.INIT_04 = 256'h0000000022320232220202022202202222202002202002232202202222023222;
defparam localram4.INIT_05 = 256'h1118765432111DCBA987111321FEDC1811111111100000000000000000000000;
defparam localram4.INIT_06 = 256'h0000BA98765432111DCBA987111321FEDC1118765432111DCBA987111321FEDC;
defparam localram4.INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;


RAMB16_S4 localram5(
	.DO     (data_out[23:20]),
	.ADDR   (addr[13:2]),
	.CLK    (clk),
	.DI     (data_in[23:20]),
	.EN     (en),
	.SSR    (reset),
	.WE     (we[2])
);
defparam localram5.INIT_00 = 256'hAAAAAAAAAAAAAA00BBBBBBBBBBBAAAAAAAAAAAAAAAB000808688B1A080910000;
defparam localram5.INIT_01 = 256'hCC040880440C060CC008804400604040CCCCABB0EBBCABB9611BBBBBBBBBBBBA;
defparam localram5.INIT_02 = 256'hC0060C400CC0048600CC4048600CCC00CCC60CCC00CC00880440C40880440040;
defparam localram5.INIT_03 = 256'h08400C8640880440C40C60C0C60CC040040C0440CC40C0060C0C40CCC040C00C;
defparam localram5.INIT_04 = 256'h00000000600608408608400C840880440C40C00C40C0460CC008804406084086;
defparam localram5.INIT_05 = 256'h0002222222000111111100011100000A00000000000000000000000000000000;
defparam localram5.INIT_06 = 256'h0000666666666600055555550005554444000444444400033333330003332222;
defparam localram5.INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;


RAMB16_S4 localram6(
	.DO     (data_out[27:24]),
	.ADDR   (addr[13:2]),
	.CLK    (clk),
	.DI     (data_in[27:24]),
	.EN     (en),
	.SSR    (reset),
	.WE     (we[3])
);
defparam localram6.INIT_00 = 256'hFFFFFFFFFFFFFF0CFFFFFFFFFFFFFFFFFFFFFFFFFF780C04440C7C4C4C7C0000;
defparam localram6.INIT_01 = 256'hFF000FF0C4CF044FF00FF0C4C044CCCCFFFF3F7037F33F703047FFFFFFFFFFFF;
defparam localram6.INIT_02 = 256'hF4040F000FF00C040CFF00C040CFFF08FFF00FFF00FF00FF0C4CF00FF0C4C000;
defparam localram6.INIT_03 = 256'h0F000FF04CFF0C4CF40FC0FCF0CFF0CC040F0480FF40F08C0FCF00FFF0CCF00F;
defparam localram6.INIT_04 = 256'h00000008C4CC0F4CF00F000FF00FF0C4CF40F08F40F0404FF00FF0C4CC0F4CF0;
defparam localram6.INIT_05 = 256'hA988765432A98DCBA987A98321FEDCA081111111100000000000000000000000;
defparam localram6.INIT_06 = 256'h0000BA98765432A98DCBA987A98321FEDCA988765432A98DCBA987A98321FEDC;
defparam localram6.INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;


RAMB16_S4 localram7(
	.DO     (data_out[31:28]),
	.ADDR   (addr[13:2]),
	.CLK    (clk),
	.DI     (data_in[31:28]),
	.EN     (en),
	.SSR    (reset),
	.WE     (we[3])
);
defparam localram7.INIT_00 = 256'h8888888888888800AAAAAAAAAAAAAAAAAAAAAAAAAA200043210A333333330101;
defparam localram7.INIT_01 = 256'h8A0308A0833A0128A008A083301283A3AAAA0A2002800A240432888888888888;
defparam localram7.INIT_02 = 256'hA201080008A00802038A30802038AA00AAA0088A008A008A0833A308A0833010;
defparam localram7.INIT_03 = 256'h080008A0338A0833A208A083A038A083010801208A20800A083A0088A083A008;
defparam localram7.INIT_04 = 256'h00000000A23A0833A0080008A308A0833A20800A20801038A008A0833A0833A0;
defparam localram7.INIT_05 = 256'h3330000000222000000011100000000C00000000000000000000000000000000;
defparam localram7.INIT_06 = 256'h0000000000000088800000007770000000666000000055500000004440000000;
defparam localram7.INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;



endmodule