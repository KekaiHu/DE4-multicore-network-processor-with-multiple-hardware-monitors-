//
// Designed by Qiang Wu
//	16K bytes, 32bit interface

`timescale 1ns/1ps


module nexthop(clk, addr, data_in, data_out, we, en, reset);
input clk;
input [13:2] addr;
input [31:0] data_in;
output [31:0] data_out;
input [3:0] we;
input en;
input reset;


RAMB16_S4 localram0(
	.DO     (data_out[3:0]),
	.ADDR   (addr[13:2]),
	.CLK    (clk),
	.DI     (data_in[3:0]),
	.EN     (en),
	.SSR    (reset),
	.WE     (we[0])
);
defparam localram0.INIT_00 = 256'h0000000000000000000000000000000000000000000000011111111111111111;
defparam localram0.INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram0.INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;


RAMB16_S4 localram1(
	.DO     (data_out[7:4]),
	.ADDR   (addr[13:2]),
	.CLK    (clk),
	.DI     (data_in[7:4]),
	.EN     (en),
	.SSR    (reset),
	.WE     (we[0])
);
defparam localram1.INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram1.INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;


RAMB16_S4 localram2(
	.DO     (data_out[11:8]),
	.ADDR   (addr[13:2]),
	.CLK    (clk),
	.DI     (data_in[11:8]),
	.EN     (en),
	.SSR    (reset),
	.WE     (we[1])
);
defparam localram2.INIT_00 = 256'h0000000000000000000000000000000000000000000000044C00C404CC488000;
defparam localram2.INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram2.INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;


RAMB16_S4 localram3(
	.DO     (data_out[15:12]),
	.ADDR   (addr[13:2]),
	.CLK    (clk),
	.DI     (data_in[15:12]),
	.EN     (en),
	.SSR    (reset),
	.WE     (we[1])
);
defparam localram3.INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram3.INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;


RAMB16_S4 localram4(
	.DO     (data_out[19:16]),
	.ADDR   (addr[13:2]),
	.CLK    (clk),
	.DI     (data_in[19:16]),
	.EN     (en),
	.SSR    (reset),
	.WE     (we[2])
);
defparam localram4.INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram4.INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;


RAMB16_S4 localram5(
	.DO     (data_out[23:20]),
	.ADDR   (addr[13:2]),
	.CLK    (clk),
	.DI     (data_in[23:20]),
	.EN     (en),
	.SSR    (reset),
	.WE     (we[2])
);
defparam localram5.INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram5.INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;


RAMB16_S4 localram6(
	.DO     (data_out[27:24]),
	.ADDR   (addr[13:2]),
	.CLK    (clk),
	.DI     (data_in[27:24]),
	.EN     (en),
	.SSR    (reset),
	.WE     (we[3])
);
defparam localram6.INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram6.INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;


RAMB16_S4 localram7(
	.DO     (data_out[31:28]),
	.ADDR   (addr[13:2]),
	.CLK    (clk),
	.DI     (data_in[31:28]),
	.EN     (en),
	.SSR    (reset),
	.WE     (we[3])
);
defparam localram7.INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam localram7.INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;



endmodule